//////////////////////////////////////////////////////////////////////////////////
// University of Toronto
// NES APU UNIT
// Engineer: Cedomir Segulja
// Create Date: 03/21/2008 
// Design Name: NES APU UNIT
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Random Generator for the Noise Channel
//////////////////////////////////////////////////////////////////////////////////

module random_generator(
                        iClk,
								iReset,
								iEnable,
								iMode,
								oData
								);
								
  //-------------------------------------------------------------------------------------------------------
  //  PORTS
  //-------------------------------------------------------------------------------------------------------

  input iClk;
  input iReset;
  input iEnable;
  input iMode;
  output oData;
  
  //-------------------------------------------------------------------------------------------------------
  //  PARAMETERS
  //-------------------------------------------------------------------------------------------------------
  
  parameter sequence_32767 = 0;
  parameter sequence_93 = 1;
  
  //-------------------------------------------------------------------------------------------------------
  //  SHIFT REGISTER
  //-------------------------------------------------------------------------------------------------------
  
  reg [14:0] shift_register;
  
  always @(posedge iClk or posedge iReset)
  begin
    if (iReset == 1)
	 begin
	   shift_register <= 15'b100000000000000;
	 end else
	 begin
	   if (iEnable)
		begin
	     if (iMode == sequence_32767)
	       shift_register[14] <= shift_register[0] ^ shift_register[1];
		  else
		    shift_register[14] <= shift_register[0] ^ shift_register[6];
		  shift_register[13:0] <= shift_register[14:1];
	   end
	 end
  end
  
  //-------------------------------------------------------------------------------------------------------
  //  OUTPUT
  //-------------------------------------------------------------------------------------------------------
  
  assign oData = !shift_register[0];

endmodule
