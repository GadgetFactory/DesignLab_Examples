//////////////////////////////////////////////////////////////////////////////////
// University of Toronto
// NES APU UNIT
// Engineer: Cedomir Segulja
// Create Date: 03/21/2008 
// Design Name: NES APU UNIT
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Trigger oChange when iSignal changes
//////////////////////////////////////////////////////////////////////////////////

module comparator(
                  iClk,
						iSignal,
						oChange
						);

  //-------------------------------------------------------------------------------------------------------
  //  PARAMETERS 
  //-------------------------------------------------------------------------------------------------------
  
  parameter WIDTH = 4;
						
  //-------------------------------------------------------------------------------------------------------
  //  PORTS
  //-------------------------------------------------------------------------------------------------------

  input iClk;
  input iSignal;
  output oChange;

  //-------------------------------------------------------------------------------------------------------
  //  REGISTERS
  //-------------------------------------------------------------------------------------------------------

  reg [WIDTH - 1:0] buffer_before;

  always @(posedge iClk)
  begin
    buffer_before <= iSignal;
  end

  //-------------------------------------------------------------------------------------------------------
  //  OUTPUT
  //-------------------------------------------------------------------------------------------------------

  assign oChange = (buffer_before == iSignal) ? 0:1;

endmodule
